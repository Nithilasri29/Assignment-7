module subtract_2s_complement (
    input  [3:0] A,
    input  [3:0] B,
    output [3:0] Result,
    output Carry
);

    wire [3:0] B_comp;
    wire [4:0] Sum;

   
    assign B_comp = ~B + 1'b1;
    assign Sum = A + B_comp;
    assign Result = Sum[3:0];
    assign Carry  = Sum[4];  

endmodule


